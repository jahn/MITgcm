netcdf grid {
dimensions:
	Z = 15 ;
	Zp1 = 16 ;
	Zu = 15 ;
	Zl = 15 ;
	X = 384 ;
	Y = 16 ;
	Xp1 = 385 ;
	Yp1 = 17 ;
variables:
	double Z(Z) ;
		Z:long_name = "vertical coordinate of cell center" ;
		Z:units = "meters" ;
		Z:positive = "up" ;
	double RC(Z) ;
		RC:description = "R coordinate of cell center" ;
		RC:units = "m" ;
	double Zp1(Zp1) ;
		Zp1:long_name = "vertical coordinate of cell interface" ;
		Zp1:units = "meters" ;
		Zp1:positive = "up" ;
	double RF(Zp1) ;
		RF:description = "R coordinate of cell interface" ;
		RF:units = "m" ;
	double Zu(Zu) ;
		Zu:long_name = "vertical coordinate of lower cell interface" ;
		Zu:units = "meters" ;
		Zu:positive = "up" ;
	double RU(Zu) ;
		RU:description = "R coordinate of upper interface" ;
		RU:units = "m" ;
	double Zl(Zl) ;
		Zl:long_name = "vertical coordinate of upper cell interface" ;
		Zl:units = "meters" ;
		Zl:positive = "up" ;
	double RL(Zl) ;
		RL:description = "R coordinate of lower interface" ;
		RL:units = "m" ;
	double drC(Zp1) ;
		drC:description = "r cell center separation" ;
	double drF(Z) ;
		drF:description = "r cell face separation" ;
	double X(X) ;
		X:long_name = "i-index of cell center" ;
		X:units = "none" ;
	double Y(Y) ;
		Y:long_name = "j-index of cell center" ;
		Y:units = "none" ;
	double XC(Y, X) ;
		XC:description = "X coordinate of cell center (T-P point)" ;
		XC:units = "degree_east" ;
	double YC(Y, X) ;
		YC:description = "Y coordinate of cell center (T-P point)" ;
		YC:units = "degree_north" ;
	double Xp1(Xp1) ;
		Xp1:long_name = "i-index of cell corner" ;
		Xp1:units = "none" ;
	double Yp1(Yp1) ;
		Yp1:long_name = "j-index of cell corner" ;
		Yp1:units = "none" ;
	double XG(Yp1, Xp1) ;
		XG:description = "X coordinate of cell corner (Vorticity point)" ;
		XG:units = "degree_east" ;
	double YG(Yp1, Xp1) ;
		YG:description = "Y coordinate of cell corner (Vorticity point)" ;
		YG:units = "degree_north" ;
	double dxC(Y, Xp1) ;
		dxC:description = "x cell center separation" ;
	double dyC(Yp1, X) ;
		dyC:description = "y cell center separation" ;
	double dxF(Y, X) ;
		dxF:description = "x cell face separation" ;
	double dyF(Y, X) ;
		dyF:description = "y cell face separation" ;
	double dxG(Yp1, X) ;
		dxG:description = "x cell corner separation" ;
	double dyG(Y, Xp1) ;
		dyG:description = "y cell corner separation" ;
	double dxV(Yp1, Xp1) ;
		dxV:description = "x v-velocity separation" ;
	double dyU(Yp1, Xp1) ;
		dyU:description = "y u-velocity separation" ;
	double rA(Y, X) ;
		rA:description = "r-face area at cell center" ;
	double rAw(Y, Xp1) ;
		rAw:description = "r-face area at U point" ;
	double rAs(Yp1, X) ;
		rAs:description = "r-face area at V point" ;
	double rAz(Yp1, Xp1) ;
		rAz:description = "r-face area at cell corner" ;
	double AngleCS(Y, X) ;
		AngleCS:description = "Cos of grid orientation angle at cell center" ;
	double AngleSN(Y, X) ;
		AngleSN:description = "Sin of grid orientation angle at cell center" ;
	double fCori(Y, X) ;
		fCori:description = "Coriolis f at cell center" ;
	double fCoriG(Yp1, Xp1) ;
		fCoriG:description = "Coriolis f at cell corner" ;
	double R_low(Y, X) ;
		R_low:description = "base of fluid in r-units" ;
	double Ro_surf(Y, X) ;
		Ro_surf:description = "surface reference (at rest) position" ;
	double Depth(Y, X) ;
		Depth:description = "fluid thickness in r coordinates (at rest)" ;
	double HFacC(Z, Y, X) ;
		HFacC:description = "vertical fraction of open cell at cell center" ;
	double HFacW(Z, Y, Xp1) ;
		HFacW:description = "vertical fraction of open cell at West face" ;
	double HFacS(Z, Yp1, X) ;
		HFacS:description = "vertical fraction of open cell at South face" ;

// global attributes:
		:MITgcm_version = "checkpoint67u" ;
		:MITgcm_URL = "http://mitgcm.org" ;
		:MITgcm_tag_id = "" ;
		:MITgcm_mnc_ver = 0.9 ;
		:sNx = 32 ;
		:sNy = 16 ;
		:OLx = 4 ;
		:OLy = 4 ;
		:nSx = 12 ;
		:nSy = 1 ;
		:nPx = 1 ;
		:nPy = 1 ;
		:Nx = 384 ;
		:Ny = 16 ;
		:Nr = 15 ;
}
