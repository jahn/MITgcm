netcdf state.0000072000 {
dimensions:
	X = 384 ;
	Y = 16 ;
	Xp1 = 385 ;
	Yp1 = 17 ;
	T = UNLIMITED ; // (2 currently)
	Z = 15 ;
	Zl = 15 ;
variables:
	double X(X) ;
		X:long_name = "i-index of cell center" ;
		X:units = "none" ;
	double Y(Y) ;
		Y:long_name = "j-index of cell center" ;
		Y:units = "none" ;
	float XC(Y, X) ;
		XC:description = "X coordinate of cell center (T-P point)" ;
		XC:units = "degree_east" ;
	float YC(Y, X) ;
		YC:description = "Y coordinate of cell center (T-P point)" ;
		YC:units = "degree_north" ;
	double Xp1(Xp1) ;
		Xp1:long_name = "i-index of cell corner" ;
		Xp1:units = "none" ;
	double Yp1(Yp1) ;
		Yp1:long_name = "j-index of cell corner" ;
		Yp1:units = "none" ;
	float XG(Yp1, Xp1) ;
		XG:description = "X coordinate of cell corner (Vorticity point)" ;
		XG:units = "degree_east" ;
	float YG(Yp1, Xp1) ;
		YG:description = "Y coordinate of cell corner (Vorticity point)" ;
		YG:units = "degree_north" ;
	double Z(Z) ;
		Z:long_name = "vertical coordinate of cell center" ;
		Z:units = "meters" ;
		Z:positive = "up" ;
	double Zl(Zl) ;
		Zl:long_name = "vertical coordinate of upper cell interface" ;
		Zl:units = "meters" ;
		Zl:positive = "up" ;
	double T(T) ;
		T:long_name = "model_time" ;
		T:units = "s" ;
	int iter(T) ;
		iter:long_name = "iteration_count" ;
	float U(T, Z, Y, Xp1) ;
		U:units = "m/s" ;
		U:coordinates = "XU YU RC iter" ;
	float V(T, Z, Yp1, X) ;
		V:units = "m/s" ;
		V:coordinates = "XV YV RC iter" ;
	float Temp(T, Z, Y, X) ;
		Temp:units = "degC" ;
		Temp:long_name = "potential_temperature" ;
		Temp:coordinates = "XC YC RC iter" ;
	float S(T, Z, Y, X) ;
		S:long_name = "salinity" ;
		S:coordinates = "XC YC RC iter" ;
	float Eta(T, Y, X) ;
		Eta:long_name = "free-surface_r-anomaly" ;
		Eta:units = "m" ;
		Eta:coordinates = "XC YC iter" ;
	float W(T, Zl, Y, X) ;
		W:units = "m/s" ;
		W:coordinates = "XC YC RC iter" ;

// global attributes:
		:MITgcm_version = "checkpoint67u" ;
		:MITgcm_URL = "http://mitgcm.org" ;
		:MITgcm_tag_id = "" ;
		:MITgcm_mnc_ver = 0.9 ;
		:sNx = 32 ;
		:sNy = 16 ;
		:OLx = 4 ;
		:OLy = 4 ;
		:nSx = 12 ;
		:nSy = 1 ;
		:nPx = 1 ;
		:nPy = 1 ;
		:Nx = 384 ;
		:Ny = 16 ;
		:Nr = 15 ;
}
